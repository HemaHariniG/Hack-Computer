module mux16_gate(a, b, sel, out);
    input [15:0] a, b;
    input sel;
    output [15:0] out;
    
    mux_gate mux0(a[0], b[0], sel, out[0]);
    mux_gate mux1(a[1], b[1], sel, out[1]);
    mux_gate mux2(a[2], b[2], sel, out[2]);
    mux_gate mux3(a[3], b[3], sel, out[3]);
    mux_gate mux4(a[4], b[4], sel, out[4]);
    mux_gate mux5(a[5], b[5], sel, out[5]);
    mux_gate mux6(a[6], b[6], sel, out[6]);
    mux_gate mux7(a[7], b[7], sel, out[7]);
    mux_gate mux8(a[8], b[8], sel, out[8]);
    mux_gate mux9(a[9], b[9], sel, out[9]);
    mux_gate mux10(a[10], b[10], sel, out[10]);
    mux_gate mux11(a[11], b[11], sel, out[11]);
    mux_gate mux12(a[12], b[12], sel, out[12]);
    mux_gate mux13(a[13], b[13], sel, out[13]);
    mux_gate mux14(a[14], b[14], sel, out[14]);
    mux_gate mux15(a[15], b[15], sel, out[15]);
endmodule
